module inststruction_mem(PC,)
input [31:0] PC;


endmodule