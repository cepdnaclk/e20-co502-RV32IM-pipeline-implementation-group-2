module imidiateGenarator(INSTRUCTION,IMMEDIATE_TYPE,IMMEDIATE_VALUE);
input [31:0] INSTRUCTION;
input [2:0] IMMEDIATE_TYPE;
output reg[31:0] IMMEDIATE_VALUE;

always @(INSTRUCTION,IMMEDIATE_TYPE) begin
    case (IMMEDIATE_TYPE)

        3'b000: IMMEDIATE_VALUE = {{21{INSTRUCTION[31]}},INSTRUCTION[30:25],INSTRUCTION[24:21],INSTRUCTION[20]};
        3'b001: IMMEDIATE_VALUE = {{21{INSTRUCTION[31]}},INSTRUCTION[30:25],INSTRUCTION[11:8],INSTRUCTION[7]};
        3'b010: IMMEDIATE_VALUE = {{12{INSTRUCTION[31]}},INSTRUCTION[19:12],INSTRUCTION[20],INSTRUCTION[30:25],INSTRUCTION[24:21],1'b0};
        3'b011: IMMEDIATE_VALUE = {INSTRUCTION[31],INSTRUCTION[30:20],INSTRUCTION[19:12],12'b0};
        3'b100: IMMEDIATE_VALUE = {{20{INSTRUCTION[31]}},INSTRUCTION[7],INSTRUCTION[30:25],INSTRUCTION[11:8],1'b0};
        
    endcase


    end


endmodule