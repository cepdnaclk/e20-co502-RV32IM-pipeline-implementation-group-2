module inststruction_mem(PC,)