module detector(PREV_INST,)